library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity seg is
port( 	BCD:in std_logic_vector(3 downto 0 );
		seg:out std_logic_vector(7 downto 0));
end seg;

architecture BCD_seg of seg is
    begin
       seg<="00000011" when bcd="0000" else
            "10011111" when bcd="0001" else
            "00100101" when bcd="0010" else
            "00001101" when bcd="0011" else
            "10011001" when bcd="0100" else
            "01001001" when bcd="0101" else
            "01000001" when bcd="0110" else
            "00011111" when bcd="0111" else
            "00000001" when bcd="1000" else
            "00001001" when bcd="1001" else
            null ;
    
end BCD_seg;