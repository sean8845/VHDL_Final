library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity t01 is
port( 	sw:in std_logic_vector(7 downto 0 );
		led:out std_logic_vector(7 downto 0));
end t01;

architecture a of t01 is
    begin
      led<=sw;
end a;